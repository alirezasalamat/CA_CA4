`timescale 1 ns / 1 ns
module datapath(clk, rst);
    input clk, rst;
    pc program_counter();

endmodule